module pratica3 (
	input wire [9:0] SW
);

contaUns();

endmodule